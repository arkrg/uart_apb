package apb_pkg;
  localparam int NUM_COMP = 5;
  localparam int ADDR_WIDTH = 32;
  localparam int DATA_WIDTH = 32;
endpackage
